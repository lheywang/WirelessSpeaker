* C:\Users\leona\Documents\.Nextcloud\Leonard\3. Projets\Enceinte\Simulations\QSPICE\schematic\top.qsch
V1 N05 0 -7
V2 N06 0 7
V3 R+ N01 AC=1 SIN 0 3.3 5000
X�Channel_SE_Filter_R+ +7V R+ -7V R+High R+Mediums R+Bass Channel_SE_Filter
X�Channel_SE_Filter_R- +7V R- -7V R-High R-Mediums R-Bass Channel_SE_Filter
X�Channel_SE_Filter_L+ +7V L+ -7V L+High L+Mediums L+Bass Channel_SE_Filter
X�Channel_SE_Filter_L- +7V L- -7V L-High L-Mediums L-Bass Channel_SE_Filter
V4 R- N01 AC=1 SIN 0 3.3 5000
V5 N01 0 {DC}
V6 L+ N02 AC=1 SIN 0 3.3 5000
V7 L- N02 AC=1 SIN 0 3.3 5000
V8 N02 0 {DC}
X�Amp_RHigh +7V -7V R+High R+High OUTR+High OUTR-High Channel_Amplifier WiperA = {wiper} WiperB = {wiper} WiperRes = {Res}
X�Amp_RMediums +7V -7V R+Mediums R-Mediums OUTR+Mediums OUTR-Mediums Channel_Amplifier WiperA = {wiper} WiperB = {wiper} WiperRes = {Res}
X�Amp_LHigh +7V -7V L+High L+High OUTL+High OUTL-High Channel_Amplifier WiperA = {wiper} WiperB = {wiper} WiperRes = {Res}
X�Amp_LMediums +7V -7V L+Mediums L-Mediums OUTL+Mediums OUTL-Mediums Channel_Amplifier WiperA ={wiper} WiperB = {wiper} WiperRes = {Res}
X�Bass_Adder +7V -7V R+Bass R-Bass N03 N04 L+Bass L-Bass Channel_Combiner
X�Amp_Bass +7V -7V N03 N04 OUT+Bass OUT-Bass Channel_Amplifier WiperA = {wiper} WiperB = {wiper} WiperRes = {Res}
V9 +7V N06 SIN 0 {AMP} 1000000
V10 -7V N05 SIN 0 {AMP} 1000000

.subckt Channel_Amplifier + - IN+ IN- OUT+ OUT-
�2 + - OUT+ N01 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
R3 N02 OUT+ (45K - {WiperA}) * {R_tol}
R4 IN+ N02 {WiperA} *  {R_tol}
�3 + - OUT- N03 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
R7 N04 OUT- (45K - {WiperB}) * {R_tol}
R8 IN- N04 {WiperB} *  {R_tol}
R1 N01 OUT+ 1.5K * {R_tol}
R2 N03 OUT- 1.5K * {R_tol}
R5 N02 N01 {WiperRes} * {R_tol}
R6 N04 N03 {WiperRes} * {R_tol}
.ends Channel_Amplifier


.subckt Channel_Combiner + - IN1+ IN1- OUT+ OUT- IN2+ IN2-
�2 + - OUT+ N01 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
�1 + - OUT- N02 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
R1 IN1+ N01 1K * {R_tol}
R2 IN2+ N01 1K * {R_tol}
R3 N01 OUT+ 2.2K * {R_tol}
R4 N02 OUT- 2.2K * {R_tol}
R5 IN2- N02 1K * {R_tol}
R6 IN1- N02 1K * {R_tol}
.ends Channel_Combiner


.subckt Channel_SE_Filter + IN - HIGH MEDIUMS BASS
X�Reconstruction_filter IN N01 + - Reconstruction_filter
X�Input_High_Pass N01 N02 + - RC_7Hz_HP
X�Bass_Filter N02 BASS + - MFB_Bass
X�Medium_Filter N02 MEDIUMS + - MFB_Mediums
X�Trebbles_Filter N02 HIGH + - MFB_High
 .subckt MFB_Bass IN OUT + -
 R3 N03 N05 470 * {R_tol}
 C3 N05 0 3.3� * {C_tol}
 �1 + - OUT N04 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C4 N01 0 820n * {C_tol}
 C5 N03 N02 100n * {C_tol}
 R5 IN N01 4.7K * {R_tol}
 R6 N01 N02 2.92K * {R_tol}
 R7 N01 N03 4.7K * {R_tol}
 �2 + - N03 N02 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 R1 N04 OUT 1.5K * {R_tol}
 R2 N05 N04 1K * {R_tol}
 C1 N01 N06 68n * {C_tol}
 R4 N06 0 22 * {R_tol}
 .ends MFB_Bass
 .subckt MFB_High IN OUT + -
 �2 + - N03 N02 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C1 N01 N02 27n * {C_tol}
 C2 IN N01 27n * {C_tol}
 C3 N01 N03 27n * {C_tol}
 R1 N02 N03 4.7K * {R_tol}
 R2 0 N01 2.2K * {R_tol}
 �1 + - N06 N05 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C4 N04 N05 33n * {C_tol}
 C5 N03 N04 33n * {C_tol}
 C6 N04 N06 33n * {C_tol}
 R3 N05 N06 4.7K * {R_tol}
 R4 0 N04 2.2K * {R_tol}
 C7 N06 N07 33n * {C_tol}
 R5 N07 0 3.3K * {R_tol}
 �3 + - OUT N07 N08 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 R6 N08 OUT 920 * {R_tol}
 R7 0 N08 8.2K * {R_tol}
 .ends MFB_High
 .subckt MFB_Mediums IN OUT + -
 �2 + - N04 N03 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C1 IN N01 680n * {C_tol}
 R1 N01 0 1.82K * {R_tol}
 C2 N01 N02 220n * {C_tol}
 R2 N02 0 1.82K * {R_tol}
 C3 N02 N03 220n * {C_tol}
 C4 N02 N04 180n * {C_tol}
 R3 N03 N04 11.5K * {R_tol}
 R4 N04 N05 300 * {R_tol}
 R5 N05 N06 1.3K * {R_tol}
 R6 N06 N07 3.3K * {R_tol}
 �1 + - N08 N07 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C5 N05 0 150n * {C_tol}
 C6 N06 0 33n * {C_tol}
 C7 N07 N08 6.8n * {C_tol}
 R7 N06 N08 1.5K * {R_tol}
 R8 N08 N09 910 * {R_tol}
 R9 N09 N10 910 * {R_tol}
 �4 + - N11 N10 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C8 N09 0 82n * {C_tol}
 C9 N10 N11 15n * {C_tol}
 R10 N09 N11 1.47K * {R_tol}
 �3 + - OUT N12 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 R11 N12 OUT 732 * {R_tol}
 R12 N11 N12 1K * {R_tol}
 .ends MFB_Mediums
 .subckt RC_7Hz_HP IN OUT + -
 �4 + - OUT N02 N01 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C1 IN N01 22u * {C_tol}
 R1 N01 0 2.2k * {R_tol}
 R2 0 N02 4.7K * {R_tol}
 R3 N02 OUT 220 *{R_tol}
 .ends RC_7Hz_HP
 .subckt Reconstruction_filter IN OUT + -
 R1 IN N01 170 * {R_tol}
 C1 N01 0 27n * {C_tol}
 C2 N02 0 3.6n * {C_tol}
 C3 N04 N03 330p * {C_tol}
 R2 N01 N02 1.85k * {R_tol}
 R3 N02 N03 4.7K * {R_tol}
 R4 N02 N04 1.85k * {R_tol}
 �4 + - N04 N03 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 C4 N05 0 3.6n * {C_tol}
 C5 OUT N06 330p * {C_tol}
 R5 N04 N05 1.5k * {R_tol}
 R6 N05 N06 3.3k * {R_tol}
 R7 N05 OUT 1.5k * {R_tol}
 �1 + - OUT N06 0 � � � � � � � � � � � RRopAmp Avol={RC4558_AVOL} GBW={RC4558_GBW} Slew={RC4558_SR} Rload=2K Phi=60
 .ends Reconstruction_filter
.ends Channel_SE_Filter

.STEP PARAM R_tol list 0.99 1 1.01
.STEP PARAM C_tol list 0.9 0.95 1.05 1.1
.PARAM RC4558_SR 2200000
.PARAM RC4558_GBW 4000000
.PARAM RC4558_AVOL 10000
.AC oct 250 1 40000
.PLOT V(R+High), V(R+Bass), V(R+Mediums)
.PLOT V(R+High) + V(R+Bass) + V(R+Mediums)
.PARAM DC 0
.PARAM AMP 0
.PARAM wiper 17000
.PARAM res 160
.end
